10
3
1
0